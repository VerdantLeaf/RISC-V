`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/17/2025 10:35:55 PM
// Design Name: 
// Module Name: cpu_core
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/// @brief RV32I core that encapsulates all components of CPU
module cpu_core #(

    WORD_SIZE = 32,
    NUM_REGS = 32,
    REG_SEL = $clog2(NUM_REGS),
    NUM_WORDS = 1024,
    ADDR_SIZE = $clog2(NUM_WORDS)

    )(
    input clk,
    input rst
    );
    // Pipeline reg flush/stall
    wire flush_ifid, flush_idex, flush_exmem, flush_memwb;
    wire stall_ifid, stall_idex, stall_exmem, stall_memwb;


    wire [ADDR_SIZE - 1 : 0] branch_target;
    wire [ADDR_SIZE - 1 : 0] pc_if, pc_id, pc_ex;
    wire [WORD_SIZE - 1 : 0] instr_if, instr_id;
    wire [WORD_SIZE - 1 : 0] data1_id, data1_ex;
    wire [WORD_SIZE - 1 : 0] data2_id, data2_ex;

    // immediates
    wire [WORD_SIZE - 1 : 0] immd_id, immd_ex;

    // rs1...
    wire [WORD_SIZE - 1 : 0] rs1_id, rs1_ex;
    wire [WORD_SIZE - 1 : 0] rs2_id, rs2_ex;
    wire [WORD_SIZE - 1 : 0] rd_id, rd_ex, rd_mem, rd_wb;


    // control signals
    // terminate in ex
    wire alu_src_id, alu_src_ex;
    wire forward_select1, forward_select2;
    wire [3:0] alu_op_id, alu_op_ex;

    // terminate in mem
    wire mem_read_id, mem_read_ex, mem_read_mem;
    wire mem_write_id, mem_write_ex, mem_write_mem;
    wire branch_id, branch_ex, branch_mem;
    wire jump_id, jump_ex, jump_mem;
    wire [1:0] data_size_id, data_size_ex, data_size_mem;
    wire data_sign_id, data_sign_ex, data_sign_mem;

    // termiante in wb
    wire mem_to_reg_id, mem_to_reg_ex, mem_to_reg_mem,  mem_to_reg_wb;
    wire reg_write_id, reg_write_ex, reg_write_mem, reg_write_wb;









    // Pipeline registers and stages
    if_stage #(

        .WORD_SIZE(WORD_SIZE),
        .NUM_WORDS(NUM_WORDS),
        .ADDR_SIZE(ADDR_SIZE)

    ) instructionfetch (
        .clk(clk),
        .rst(rst),
        
        .pc_src(pc_src),
        .en(en_pc_reg), // Enables updating of PC register. Sourced from branch unit?
        
        .branch_target(branch_target),
        .pc_next(pc_if),

        .instr(instr_if)
    );

    if_id_reg #(
       
        .WORD_SIZE(WORD_SIZE)

    ) IFID_register (
        .clk(clk),
        .rst(rst),
        .flush(flush_ifid),
        .stall(stall_ifid),

        .instr(instr_if),
        .pc(pc_if),

        .instr_out(instr_id), // instruction and PC to ID stage
        .pc_out(pc_id)
    );

    id_stage #(
        .WORD_SIZE(WORD_SIZE),
        .NUM_REGS(NUM_REGS),
        .NUM_WORDS(NUM_WORDS),
        .REG_SEL(REG_SEL),
        .ADDR_SIZE(ADDR_SIZE)
    ) instructiondecode (
        .clk(clk),
        .rst(rst),

        .instr(instr_id),

        .reg_write(),
        .rd_data(),
        .rd_select(rd_wb),

        .immd(immd_id),
        .data1(),
        .data2(),
        .alu_op(alu_op_id),
        .rd(rd_id),
        .rs1(rs1_id),
        .rs2(rs2_id),

        .mem_read(mem_read_id),
        .mem_write(mem_write_id),
        .mem_to_reg(mem_to_reg_id),
        .reg_write(reg_write_id),
        .alu_src(alu_src_id),
        .branch(branch_id),
        .jump(jump_id),

        .data_size(data_size_id),
        .data_sign(data_sign_id),
    );

    id_ex_reg #(

        .WORD_SIZE(WORD_SIZE),
        .NUM_REGS(NUM_REGS),
        .NUM_WORDS(NUM_WORDS),
        .REG_SEL(NUM_REGS),
        .ADDR_SIZE(ADDR_SIZE)

    ) IDEX_register (
        .clk(clk),
        .rst(rst),
        .flush(flush_idex),
        .stall(stall_idex),

        .pc(pc_id),
        .immd(immd_id),
        .data1(),
        .data2(),

        .alu_op(alu_op_id),
        .rd(rd_id),
        .rs1(rs1_id),
        .rs2(rs2_id),

        .mem_read(mem_read_id),
        .mem_write(mem_write_id),
        .mem_to_reg(mem_to_reg_id),
        .reg_write(reg_write_id),
        .alu_src(alu_src_id),
        .branch(branch_id),
        .jump(jump_id),

        .data_size(data_size_id),
        .data_sign(data_sign_id),

        .pc_out(pc_ex),
        .immd_out(),
        .data1_out(),
        .data2_out(),

        .alu_op_out(alu_op_ex),
        .rs1_out(rs1_ex),
        .rs2_out(rs2_ex),
        .rd_out(rd_ex),

        .mem_read_out(mem_read_ex),
        .mem_write_out(mem_write_ex),
        .mem_to_reg_out(mem_to_reg_ex),
        .reg_write_out(reg_write_ex),
        .alu_src_out(alu_src_ex),
        .branch_out(branch_ex),
        .jump_out(jump_ex),
        
        .data_size_out(data_size_ex),
        .data_sign_out(data_sign_ex)

    );

    ex_stage #(
        .WORD_SIZE(WORD_SIZE),
        .NUM_REGS(NUM_REGS),
        .NUM_WORDS(NUM_WORDS),
        .REG_SEL(NUM_REGS),
        .ADDR_SIZE(ADDR_SIZE)
    )execution(
        .pc(pc_ex),
    );

    ex_mem_reg #(
        .WORD_SIZE(WORD_SIZE),
        .NUM_REGS(NUM_REGS),
        .NUM_WORDS(NUM_WORDS),
        .REG_SEL(REG_SEL),
        .ADDR_SIZE(ADDR_SIZE)
    ) EXMEM_register (
        .clk(clk),
        .rst(rst),
        .flush(flush_exmem),
        .stall(stall_exmem),

        .branch_target(),
        .alu_result(),
        .rd(rd_ex),

        .mem_read(),
        .mem_write(),
        .mem_to_reg(),
        .reg_write(),
        .alu_zero(),
        .branch(),
        .jump(),

        .write_data(),
        .data_size(data_size_ex),
        .data_sign(data_sign_ex),


        .branch_target_out(),
        .alu_result_out(),
        .rd_out(rd_mem),

        .mem_read_out(),
        .mem_write_out(),
        .mem_to_reg_out(),
        .reg_write_out(),
        .alu_zero_out(),
        .branch_out(),
        .jump_out(),

        .write_data_out(),
        .data_size_out(data_size_mem),
        .data_sign_out(data_sign_mem)
    );

    mem_stage memory();

    mem_wb_reg #(

    ) MEMWB_register (
        
        .rd(rd_mem),

        .rd(rd_wb)
    );

    wb_stage #(
        .WORD_SIZE(WORD_SIZE)
    )writeback(
        .memory_data(read_data),
        .alu_data(alu_res_wb),
        .mem_to_reg(mem_to_reg_wb),
        .write_data(write_data_to_regfile)
    );

    // External control and hazard units
    forwarding_unit forwarding_unit();

    branch_unit branch_unit();

endmodule
